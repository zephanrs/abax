module __mv__mv_0_next(
  input wire clk,
  input wire rst,
  input wire mv__done_rdy,
  input wire mv__go,
  input wire mv__go_vld,
  input wire mv__mem0__read_req_rdy,
  input wire [31:0] mv__mem0__read_resp,
  input wire mv__mem0__read_resp_vld,
  input wire mv__mem1__read_req_rdy,
  input wire [31:0] mv__mem1__read_resp,
  input wire mv__mem1__read_resp_vld,
  input wire mv__mem2__write_req_rdy,
  input wire mv__mem2__write_resp_vld,
  output wire mv__done,
  output wire mv__done_vld,
  output wire mv__go_rdy,
  output wire [3:0] mv__mem0__read_req,
  output wire mv__mem0__read_req_vld,
  output wire mv__mem0__read_resp_rdy,
  output wire [1:0] mv__mem1__read_req,
  output wire mv__mem1__read_req_vld,
  output wire mv__mem1__read_resp_rdy,
  output wire [33:0] mv__mem2__write_req,
  output wire mv__mem2__write_req_vld,
  output wire mv__mem2__write_resp_rdy
);
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [31:0] smul32b_32b_x_32b (input reg [31:0] lhs, input reg [31:0] rhs);
    reg signed [31:0] signed_lhs;
    reg signed [31:0] signed_rhs;
    reg signed [31:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul32b_32b_x_32b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  wire [31:0] __mv__mem0__read_resp_reg_init = 32'h0000_0000;
  wire [31:0] __mv__mem1__read_resp_reg_init = 32'h0000_0000;
  wire [3:0] __mv__mem0__read_req_reg_init = 4'h0;
  wire [1:0] __mv__mem1__read_req_reg_init = 2'h0;
  wire [33:0] __mv__mem2__write_req_reg_init = {2'h0, 32'h0000_0000};
  reg [31:0] ____state_1;
  reg [1:0] ____state_2;
  reg ____state_3;
  reg [1:0] p0_tmp21;
  reg p0_or_534;
  reg p0_and_552;
  reg p0_tmp25;
  reg p0_and_546;
  reg [1:0] p1_tmp21;
  reg p1_or_534;
  reg [31:0] p1_tmp15;
  reg p1_and_552;
  reg p1_tmp25;
  reg p1_and_546;
  reg [31:0] ____state_0;
  reg p2_and_552;
  reg p2_tmp25;
  reg p0_valid;
  reg p1_valid;
  reg p2_valid;
  reg __mv__mem0__read_req_has_been_sent_reg;
  reg __mv__mem1__read_req_has_been_sent_reg;
  reg __mv__mem2__write_req_has_been_sent_reg;
  reg __mv__done_has_been_sent_reg;
  reg __mv__go_reg;
  reg __mv__go_valid_reg;
  reg [31:0] __mv__mem0__read_resp_reg;
  reg __mv__mem0__read_resp_valid_reg;
  reg [31:0] __mv__mem1__read_resp_reg;
  reg __mv__mem1__read_resp_valid_reg;
  reg __mv__mem2__write_resp_valid_reg;
  reg [3:0] __mv__mem0__read_req_reg;
  reg __mv__mem0__read_req_valid_reg;
  reg [1:0] __mv__mem1__read_req_reg;
  reg __mv__mem1__read_req_valid_reg;
  reg [33:0] __mv__mem2__write_req_reg;
  reg __mv__mem2__write_req_valid_reg;
  reg __mv__done_reg;
  reg __mv__done_valid_reg;
  wire or_650;
  wire __mv__done_vld_buf;
  wire __mv__done_not_has_been_sent;
  wire mv__done_valid_inv;
  wire __mv__done_valid_and_not_has_been_sent;
  wire mv__done_valid_load_en;
  wire mv__done_load_en;
  wire or_879;
  wire p3_stage_done;
  wire p3_not_valid;
  wire p2_enable;
  wire __mv__mem2__write_req_vld_buf;
  wire __mv__mem2__write_req_not_has_been_sent;
  wire mv__mem2__write_req_valid_inv;
  wire __mv__mem2__write_req_valid_and_not_has_been_sent;
  wire mv__mem2__write_req_valid_load_en;
  wire mv__mem2__write_req_load_en;
  wire or_878;
  wire p2_stage_done;
  wire p2_data_enable;
  wire p2_not_valid;
  wire p1_all_active_inputs_valid;
  wire p1_enable;
  wire p1_stage_done;
  wire p1_data_enable;
  wire p1_not_valid;
  wire or_646;
  wire p0_enable;
  wire __mv__mem0__read_req_vld_buf;
  wire __mv__mem0__read_req_not_has_been_sent;
  wire mv__mem0__read_req_valid_inv;
  wire __mv__mem1__read_req_not_has_been_sent;
  wire mv__mem1__read_req_valid_inv;
  wire [2:0] add_531;
  wire [31:0] add_532;
  wire __mv__mem0__read_req_valid_and_not_has_been_sent;
  wire mv__mem0__read_req_valid_load_en;
  wire __mv__mem1__read_req_valid_and_not_has_been_sent;
  wire mv__mem1__read_req_valid_load_en;
  wire tmp20;
  wire sge_536;
  wire mv__mem0__read_req_load_en;
  wire mv__mem1__read_req_load_en;
  wire nand_538;
  wire slt_539;
  wire __mv__mem0__read_req_has_sent_or_is_ready;
  wire __mv__mem1__read_req_has_sent_or_is_ready;
  wire tmp25;
  wire and_546;
  wire nor_547;
  wire p0_all_active_outputs_ready;
  wire [1:0] ____state_0__next_value_predicates;
  wire [1:0] ____state_1__next_value_predicates;
  wire [1:0] ____state_2__next_value_predicates;
  wire p0_stage_done;
  wire [2:0] one_hot_554;
  wire [2:0] one_hot_555;
  wire [2:0] one_hot_556;
  wire p0_data_enable;
  wire mv__go_select;
  wire mv__go_valid_inv;
  wire mv__mem0__read_resp_valid_inv;
  wire mv__mem1__read_resp_valid_inv;
  wire mv__mem2__write_resp_valid_inv;
  wire and_706;
  wire and_707;
  wire [31:0] tmp3;
  wire and_713;
  wire and_714;
  wire and_721;
  wire and_722;
  wire [1:0] tmp21;
  wire mv__go_valid_load_en;
  wire mv__mem0__read_resp_valid_load_en;
  wire mv__mem1__read_resp_valid_load_en;
  wire mv__mem2__write_resp_valid_load_en;
  wire ____state_0__at_most_one_next_value;
  wire ____state_1__at_most_one_next_value;
  wire ____state_2__at_most_one_next_value;
  wire [31:0] tmp6_data;
  wire [31:0] tmp10_data;
  wire [1:0] concat_709;
  wire [31:0] tmp17;
  wire [31:0] tmp2;
  wire [1:0] concat_716;
  wire tmp1;
  wire [1:0] concat_723;
  wire [1:0] unexpand_for_next_value_129_2_case_1;
  wire [1:0] unexpand_for_next_value_129_2_case_0;
  wire __mv__mem0__read_req_valid_and_all_active_outputs_ready;
  wire __mv__mem0__read_req_valid_and_ready_txfr;
  wire __mv__mem1__read_req_valid_and_ready_txfr;
  wire __mv__mem2__write_req_valid_and_all_active_outputs_ready;
  wire __mv__mem2__write_req_valid_and_ready_txfr;
  wire __mv__done_valid_and_all_active_outputs_ready;
  wire __mv__done_valid_and_ready_txfr;
  wire [3:0] tmp4;
  wire mv__go_load_en;
  wire mv__mem0__read_resp_load_en;
  wire mv__mem1__read_resp_load_en;
  wire mv__mem2__write_resp_load_en;
  wire or_873;
  wire or_875;
  wire or_877;
  wire [31:0] tmp15;
  wire or_534;
  wire and_552;
  wire [31:0] one_hot_sel_710;
  wire or_711;
  wire [31:0] one_hot_sel_717;
  wire or_718;
  wire tmp29;
  wire [1:0] one_hot_sel_724;
  wire or_725;
  wire __mv__mem0__read_req_not_stage_load;
  wire __mv__mem0__read_req_has_been_sent_reg_load_en;
  wire __mv__mem1__read_req_has_been_sent_reg_load_en;
  wire __mv__mem2__write_req_not_stage_load;
  wire __mv__mem2__write_req_has_been_sent_reg_load_en;
  wire __mv__done_not_stage_load;
  wire __mv__done_has_been_sent_reg_load_en;
  wire [3:0] tmp5;
  wire [1:0] tmp9;
  wire [33:0] tmp23;
  wire __mv__done_buf;
  assign or_650 = ~p2_and_552 | __mv__mem2__write_resp_valid_reg;
  assign __mv__done_vld_buf = or_650 & p2_valid & p2_tmp25;
  assign __mv__done_not_has_been_sent = ~__mv__done_has_been_sent_reg;
  assign mv__done_valid_inv = ~__mv__done_valid_reg;
  assign __mv__done_valid_and_not_has_been_sent = __mv__done_vld_buf & __mv__done_not_has_been_sent;
  assign mv__done_valid_load_en = mv__done_rdy | mv__done_valid_inv;
  assign mv__done_load_en = __mv__done_valid_and_not_has_been_sent & mv__done_valid_load_en;
  assign or_879 = ~p2_tmp25 | mv__done_load_en | __mv__done_has_been_sent_reg;
  assign p3_stage_done = p2_valid & or_650 & or_879;
  assign p3_not_valid = ~p2_valid;
  assign p2_enable = p3_stage_done | p3_not_valid;
  assign __mv__mem2__write_req_vld_buf = p1_valid & p2_enable & p1_and_552;
  assign __mv__mem2__write_req_not_has_been_sent = ~__mv__mem2__write_req_has_been_sent_reg;
  assign mv__mem2__write_req_valid_inv = ~__mv__mem2__write_req_valid_reg;
  assign __mv__mem2__write_req_valid_and_not_has_been_sent = __mv__mem2__write_req_vld_buf & __mv__mem2__write_req_not_has_been_sent;
  assign mv__mem2__write_req_valid_load_en = mv__mem2__write_req_rdy | mv__mem2__write_req_valid_inv;
  assign mv__mem2__write_req_load_en = __mv__mem2__write_req_valid_and_not_has_been_sent & mv__mem2__write_req_valid_load_en;
  assign or_878 = ~p1_and_552 | mv__mem2__write_req_load_en | __mv__mem2__write_req_has_been_sent_reg;
  assign p2_stage_done = p1_valid & or_878;
  assign p2_data_enable = p2_enable & p2_stage_done;
  assign p2_not_valid = ~p1_valid;
  assign p1_all_active_inputs_valid = __mv__mem0__read_resp_valid_reg & __mv__mem1__read_resp_valid_reg;
  assign p1_enable = p2_data_enable | p2_not_valid;
  assign p1_stage_done = p0_valid & p1_all_active_inputs_valid;
  assign p1_data_enable = p1_enable & p1_stage_done;
  assign p1_not_valid = ~p0_valid;
  assign or_646 = ____state_3 | __mv__go_valid_reg;
  assign p0_enable = p1_data_enable | p1_not_valid;
  assign __mv__mem0__read_req_vld_buf = or_646 & p0_enable;
  assign __mv__mem0__read_req_not_has_been_sent = ~__mv__mem0__read_req_has_been_sent_reg;
  assign mv__mem0__read_req_valid_inv = ~__mv__mem0__read_req_valid_reg;
  assign __mv__mem1__read_req_not_has_been_sent = ~__mv__mem1__read_req_has_been_sent_reg;
  assign mv__mem1__read_req_valid_inv = ~__mv__mem1__read_req_valid_reg;
  assign add_531 = {1'h0, ____state_2} + 3'h1;
  assign add_532 = ____state_1 + 32'h0000_0001;
  assign __mv__mem0__read_req_valid_and_not_has_been_sent = __mv__mem0__read_req_vld_buf & __mv__mem0__read_req_not_has_been_sent;
  assign mv__mem0__read_req_valid_load_en = mv__mem0__read_req_rdy | mv__mem0__read_req_valid_inv;
  assign __mv__mem1__read_req_valid_and_not_has_been_sent = __mv__mem0__read_req_vld_buf & __mv__mem1__read_req_not_has_been_sent;
  assign mv__mem1__read_req_valid_load_en = mv__mem1__read_req_rdy | mv__mem1__read_req_valid_inv;
  assign tmp20 = add_531[2];
  assign sge_536 = $signed(add_532) >= $signed(32'h0000_0004);
  assign mv__mem0__read_req_load_en = __mv__mem0__read_req_valid_and_not_has_been_sent & mv__mem0__read_req_valid_load_en;
  assign mv__mem1__read_req_load_en = __mv__mem1__read_req_valid_and_not_has_been_sent & mv__mem1__read_req_valid_load_en;
  assign nand_538 = ~(tmp20 & sge_536);
  assign slt_539 = $signed(____state_1) < $signed(32'h0000_0004);
  assign __mv__mem0__read_req_has_sent_or_is_ready = mv__mem0__read_req_load_en | __mv__mem0__read_req_has_been_sent_reg;
  assign __mv__mem1__read_req_has_sent_or_is_ready = mv__mem1__read_req_load_en | __mv__mem1__read_req_has_been_sent_reg;
  assign tmp25 = tmp20 & sge_536;
  assign and_546 = nand_538 & slt_539;
  assign nor_547 = ~(~tmp20 | sge_536);
  assign p0_all_active_outputs_ready = __mv__mem0__read_req_has_sent_or_is_ready & __mv__mem1__read_req_has_sent_or_is_ready;
  assign ____state_0__next_value_predicates = {tmp25, and_546};
  assign ____state_1__next_value_predicates = {tmp25, nor_547};
  assign ____state_2__next_value_predicates = {~tmp20, tmp20};
  assign p0_stage_done = or_646 & p0_all_active_outputs_ready;
  assign one_hot_554 = {____state_0__next_value_predicates[1:0] == 2'h0, ____state_0__next_value_predicates[1] && !____state_0__next_value_predicates[0], ____state_0__next_value_predicates[0]};
  assign one_hot_555 = {____state_1__next_value_predicates[1:0] == 2'h0, ____state_1__next_value_predicates[1] && !____state_1__next_value_predicates[0], ____state_1__next_value_predicates[0]};
  assign one_hot_556 = {____state_2__next_value_predicates[1:0] == 2'h0, ____state_2__next_value_predicates[1] && !____state_2__next_value_predicates[0], ____state_2__next_value_predicates[0]};
  assign p0_data_enable = p0_enable & p0_stage_done;
  assign mv__go_select = ~____state_3 ? __mv__go_reg : 1'h0;
  assign mv__go_valid_inv = ~__mv__go_valid_reg;
  assign mv__mem0__read_resp_valid_inv = ~__mv__mem0__read_resp_valid_reg;
  assign mv__mem1__read_resp_valid_inv = ~__mv__mem1__read_resp_valid_reg;
  assign mv__mem2__write_resp_valid_inv = ~__mv__mem2__write_resp_valid_reg;
  assign and_706 = p1_tmp25 & p2_data_enable;
  assign and_707 = p1_and_546 & p2_data_enable;
  assign tmp3 = ____state_0 & {32{p1_or_534}};
  assign and_713 = tmp25 & p0_data_enable;
  assign and_714 = nor_547 & p0_data_enable;
  assign and_721 = ~tmp20 & p0_data_enable;
  assign and_722 = tmp20 & p0_data_enable;
  assign tmp21 = ____state_1[1:0];
  assign mv__go_valid_load_en = p0_data_enable & ~____state_3 | mv__go_valid_inv;
  assign mv__mem0__read_resp_valid_load_en = p1_data_enable | mv__mem0__read_resp_valid_inv;
  assign mv__mem1__read_resp_valid_load_en = p1_data_enable | mv__mem1__read_resp_valid_inv;
  assign mv__mem2__write_resp_valid_load_en = p3_stage_done & p2_and_552 | mv__mem2__write_resp_valid_inv;
  assign ____state_0__at_most_one_next_value = tmp25 == one_hot_554[1] & and_546 == one_hot_554[0];
  assign ____state_1__at_most_one_next_value = tmp25 == one_hot_555[1] & nor_547 == one_hot_555[0];
  assign ____state_2__at_most_one_next_value = ~tmp20 == one_hot_556[1] & tmp20 == one_hot_556[0];
  assign tmp6_data = __mv__mem0__read_resp_reg[31:0];
  assign tmp10_data = __mv__mem1__read_resp_reg[31:0];
  assign concat_709 = {and_706, and_707};
  assign tmp17 = tmp3 + p1_tmp15;
  assign tmp2 = 32'h0000_0000;
  assign concat_716 = {and_713, and_714};
  assign tmp1 = ~(____state_3 | ~mv__go_select);
  assign concat_723 = {and_721, and_722};
  assign unexpand_for_next_value_129_2_case_1 = 2'h0;
  assign unexpand_for_next_value_129_2_case_0 = add_531[1:0];
  assign __mv__mem0__read_req_valid_and_all_active_outputs_ready = __mv__mem0__read_req_vld_buf & p0_all_active_outputs_ready;
  assign __mv__mem0__read_req_valid_and_ready_txfr = __mv__mem0__read_req_valid_and_not_has_been_sent & mv__mem0__read_req_load_en;
  assign __mv__mem1__read_req_valid_and_ready_txfr = __mv__mem1__read_req_valid_and_not_has_been_sent & mv__mem1__read_req_load_en;
  assign __mv__mem2__write_req_valid_and_all_active_outputs_ready = __mv__mem2__write_req_vld_buf & or_878;
  assign __mv__mem2__write_req_valid_and_ready_txfr = __mv__mem2__write_req_valid_and_not_has_been_sent & mv__mem2__write_req_load_en;
  assign __mv__done_valid_and_all_active_outputs_ready = __mv__done_vld_buf & or_879;
  assign __mv__done_valid_and_ready_txfr = __mv__done_valid_and_not_has_been_sent & mv__done_load_en;
  assign tmp4 = {tmp21, ____state_2};
  assign mv__go_load_en = mv__go_vld & mv__go_valid_load_en;
  assign mv__mem0__read_resp_load_en = mv__mem0__read_resp_vld & mv__mem0__read_resp_valid_load_en;
  assign mv__mem1__read_resp_load_en = mv__mem1__read_resp_vld & mv__mem1__read_resp_valid_load_en;
  assign mv__mem2__write_resp_load_en = mv__mem2__write_resp_vld & mv__mem2__write_resp_valid_load_en;
  assign or_873 = ~p0_stage_done | ____state_0__at_most_one_next_value | rst;
  assign or_875 = ~p0_stage_done | ____state_1__at_most_one_next_value | rst;
  assign or_877 = ~p0_stage_done | ____state_2__at_most_one_next_value | rst;
  assign tmp15 = smul32b_32b_x_32b(tmp6_data, tmp10_data);
  assign or_534 = ____state_2[0] | ____state_2[1];
  assign and_552 = tmp20 & slt_539;
  assign one_hot_sel_710 = tmp17 & {32{concat_709[0]}} | tmp2 & {32{concat_709[1]}};
  assign or_711 = and_706 | and_707;
  assign one_hot_sel_717 = add_532 & {32{concat_716[0]}} | tmp2 & {32{concat_716[1]}};
  assign or_718 = and_713 | and_714;
  assign tmp29 = tmp1 | ____state_3 & nand_538;
  assign one_hot_sel_724 = unexpand_for_next_value_129_2_case_1 & {2{concat_723[0]}} | unexpand_for_next_value_129_2_case_0 & {2{concat_723[1]}};
  assign or_725 = and_721 | and_722;
  assign __mv__mem0__read_req_not_stage_load = ~__mv__mem0__read_req_valid_and_all_active_outputs_ready;
  assign __mv__mem0__read_req_has_been_sent_reg_load_en = __mv__mem0__read_req_valid_and_ready_txfr | __mv__mem0__read_req_valid_and_all_active_outputs_ready;
  assign __mv__mem1__read_req_has_been_sent_reg_load_en = __mv__mem1__read_req_valid_and_ready_txfr | __mv__mem0__read_req_valid_and_all_active_outputs_ready;
  assign __mv__mem2__write_req_not_stage_load = ~__mv__mem2__write_req_valid_and_all_active_outputs_ready;
  assign __mv__mem2__write_req_has_been_sent_reg_load_en = __mv__mem2__write_req_valid_and_ready_txfr | __mv__mem2__write_req_valid_and_all_active_outputs_ready;
  assign __mv__done_not_stage_load = ~__mv__done_valid_and_all_active_outputs_ready;
  assign __mv__done_has_been_sent_reg_load_en = __mv__done_valid_and_ready_txfr | __mv__done_valid_and_all_active_outputs_ready;
  assign tmp5 = {tmp4};
  assign tmp9 = {____state_2};
  assign tmp23 = {p1_tmp21, tmp17};
  assign __mv__done_buf = 1'h1;
  always_ff @ (posedge clk) begin
    if (rst) begin
      ____state_1 <= 32'h0000_0000;
      ____state_2 <= 2'h0;
      ____state_3 <= 1'h0;
      p0_tmp21 <= 2'h0;
      p0_or_534 <= 1'h0;
      p0_and_552 <= 1'h0;
      p0_tmp25 <= 1'h0;
      p0_and_546 <= 1'h0;
      p1_tmp21 <= 2'h0;
      p1_or_534 <= 1'h0;
      p1_tmp15 <= 32'h0000_0000;
      p1_and_552 <= 1'h0;
      p1_tmp25 <= 1'h0;
      p1_and_546 <= 1'h0;
      ____state_0 <= 32'h0000_0000;
      p2_and_552 <= 1'h0;
      p2_tmp25 <= 1'h0;
      p0_valid <= 1'h0;
      p1_valid <= 1'h0;
      p2_valid <= 1'h0;
      __mv__mem0__read_req_has_been_sent_reg <= 1'h0;
      __mv__mem1__read_req_has_been_sent_reg <= 1'h0;
      __mv__mem2__write_req_has_been_sent_reg <= 1'h0;
      __mv__done_has_been_sent_reg <= 1'h0;
      __mv__go_reg <= 1'h0;
      __mv__go_valid_reg <= 1'h0;
      __mv__mem0__read_resp_reg <= __mv__mem0__read_resp_reg_init;
      __mv__mem0__read_resp_valid_reg <= 1'h0;
      __mv__mem1__read_resp_reg <= __mv__mem1__read_resp_reg_init;
      __mv__mem1__read_resp_valid_reg <= 1'h0;
      __mv__mem2__write_resp_valid_reg <= 1'h0;
      __mv__mem0__read_req_reg <= __mv__mem0__read_req_reg_init;
      __mv__mem0__read_req_valid_reg <= 1'h0;
      __mv__mem1__read_req_reg <= __mv__mem1__read_req_reg_init;
      __mv__mem1__read_req_valid_reg <= 1'h0;
      __mv__mem2__write_req_reg <= __mv__mem2__write_req_reg_init;
      __mv__mem2__write_req_valid_reg <= 1'h0;
      __mv__done_reg <= 1'h0;
      __mv__done_valid_reg <= 1'h0;
    end else begin
      ____state_1 <= or_718 ? one_hot_sel_717 : ____state_1;
      ____state_2 <= or_725 ? one_hot_sel_724 : ____state_2;
      ____state_3 <= p0_data_enable ? tmp29 : ____state_3;
      p0_tmp21 <= p0_data_enable ? tmp21 : p0_tmp21;
      p0_or_534 <= p0_data_enable ? or_534 : p0_or_534;
      p0_and_552 <= p0_data_enable ? and_552 : p0_and_552;
      p0_tmp25 <= p0_data_enable ? tmp25 : p0_tmp25;
      p0_and_546 <= p0_data_enable ? and_546 : p0_and_546;
      p1_tmp21 <= p1_data_enable ? p0_tmp21 : p1_tmp21;
      p1_or_534 <= p1_data_enable ? p0_or_534 : p1_or_534;
      p1_tmp15 <= p1_data_enable ? tmp15 : p1_tmp15;
      p1_and_552 <= p1_data_enable ? p0_and_552 : p1_and_552;
      p1_tmp25 <= p1_data_enable ? p0_tmp25 : p1_tmp25;
      p1_and_546 <= p1_data_enable ? p0_and_546 : p1_and_546;
      ____state_0 <= or_711 ? one_hot_sel_710 : ____state_0;
      p2_and_552 <= p2_data_enable ? p1_and_552 : p2_and_552;
      p2_tmp25 <= p2_data_enable ? p1_tmp25 : p2_tmp25;
      p0_valid <= p0_enable ? p0_stage_done : p0_valid;
      p1_valid <= p1_enable ? p1_stage_done : p1_valid;
      p2_valid <= p2_enable ? p2_stage_done : p2_valid;
      __mv__mem0__read_req_has_been_sent_reg <= __mv__mem0__read_req_has_been_sent_reg_load_en ? __mv__mem0__read_req_not_stage_load : __mv__mem0__read_req_has_been_sent_reg;
      __mv__mem1__read_req_has_been_sent_reg <= __mv__mem1__read_req_has_been_sent_reg_load_en ? __mv__mem0__read_req_not_stage_load : __mv__mem1__read_req_has_been_sent_reg;
      __mv__mem2__write_req_has_been_sent_reg <= __mv__mem2__write_req_has_been_sent_reg_load_en ? __mv__mem2__write_req_not_stage_load : __mv__mem2__write_req_has_been_sent_reg;
      __mv__done_has_been_sent_reg <= __mv__done_has_been_sent_reg_load_en ? __mv__done_not_stage_load : __mv__done_has_been_sent_reg;
      __mv__go_reg <= mv__go_load_en ? mv__go : __mv__go_reg;
      __mv__go_valid_reg <= mv__go_valid_load_en ? mv__go_vld : __mv__go_valid_reg;
      __mv__mem0__read_resp_reg <= mv__mem0__read_resp_load_en ? mv__mem0__read_resp : __mv__mem0__read_resp_reg;
      __mv__mem0__read_resp_valid_reg <= mv__mem0__read_resp_valid_load_en ? mv__mem0__read_resp_vld : __mv__mem0__read_resp_valid_reg;
      __mv__mem1__read_resp_reg <= mv__mem1__read_resp_load_en ? mv__mem1__read_resp : __mv__mem1__read_resp_reg;
      __mv__mem1__read_resp_valid_reg <= mv__mem1__read_resp_valid_load_en ? mv__mem1__read_resp_vld : __mv__mem1__read_resp_valid_reg;
      __mv__mem2__write_resp_valid_reg <= mv__mem2__write_resp_valid_load_en ? mv__mem2__write_resp_vld : __mv__mem2__write_resp_valid_reg;
      __mv__mem0__read_req_reg <= mv__mem0__read_req_load_en ? tmp5 : __mv__mem0__read_req_reg;
      __mv__mem0__read_req_valid_reg <= mv__mem0__read_req_valid_load_en ? __mv__mem0__read_req_valid_and_not_has_been_sent : __mv__mem0__read_req_valid_reg;
      __mv__mem1__read_req_reg <= mv__mem1__read_req_load_en ? tmp9 : __mv__mem1__read_req_reg;
      __mv__mem1__read_req_valid_reg <= mv__mem1__read_req_valid_load_en ? __mv__mem1__read_req_valid_and_not_has_been_sent : __mv__mem1__read_req_valid_reg;
      __mv__mem2__write_req_reg <= mv__mem2__write_req_load_en ? tmp23 : __mv__mem2__write_req_reg;
      __mv__mem2__write_req_valid_reg <= mv__mem2__write_req_valid_load_en ? __mv__mem2__write_req_valid_and_not_has_been_sent : __mv__mem2__write_req_valid_reg;
      __mv__done_reg <= mv__done_load_en ? __mv__done_buf : __mv__done_reg;
      __mv__done_valid_reg <= mv__done_valid_load_en ? __mv__done_valid_and_not_has_been_sent : __mv__done_valid_reg;
    end
  end
  assign mv__done = __mv__done_reg;
  assign mv__done_vld = __mv__done_valid_reg;
  assign mv__go_rdy = mv__go_load_en;
  assign mv__mem0__read_req = __mv__mem0__read_req_reg;
  assign mv__mem0__read_req_vld = __mv__mem0__read_req_valid_reg;
  assign mv__mem0__read_resp_rdy = mv__mem0__read_resp_load_en;
  assign mv__mem1__read_req = __mv__mem1__read_req_reg;
  assign mv__mem1__read_req_vld = __mv__mem1__read_req_valid_reg;
  assign mv__mem1__read_resp_rdy = mv__mem1__read_resp_load_en;
  assign mv__mem2__write_req = __mv__mem2__write_req_reg;
  assign mv__mem2__write_req_vld = __mv__mem2__write_req_valid_reg;
  assign mv__mem2__write_resp_rdy = mv__mem2__write_resp_load_en;
  `ifdef ASSERT_ON
  ____state_0__at_most_one_next_value_assert: assert property (@(posedge clk) disable iff ($sampled(rst !== 1'h0 || $isunknown(or_873))) or_873) else $fatal(0, "More than one next_value fired for state element: __state_0");
  ____state_1__at_most_one_next_value_assert: assert property (@(posedge clk) disable iff ($sampled(rst !== 1'h0 || $isunknown(or_875))) or_875) else $fatal(0, "More than one next_value fired for state element: __state_1");
  ____state_2__at_most_one_next_value_assert: assert property (@(posedge clk) disable iff ($sampled(rst !== 1'h0 || $isunknown(or_877))) or_877) else $fatal(0, "More than one next_value fired for state element: __state_2");
  `endif  // ASSERT_ON
endmodule
