module __dslx__mm4(
  input wire clk,
  input wire [511:0] a,
  input wire [511:0] b,
  output wire [511:0] out
);
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [31:0] smul32b_32b_x_32b (input reg [31:0] lhs, input reg [31:0] rhs);
    reg signed [31:0] signed_lhs;
    reg signed [31:0] signed_rhs;
    reg signed [31:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul32b_32b_x_32b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  wire [31:0] a_unflattened[4][4];
  assign a_unflattened[0][0] = a[31:0];
  assign a_unflattened[0][1] = a[63:32];
  assign a_unflattened[0][2] = a[95:64];
  assign a_unflattened[0][3] = a[127:96];
  assign a_unflattened[1][0] = a[159:128];
  assign a_unflattened[1][1] = a[191:160];
  assign a_unflattened[1][2] = a[223:192];
  assign a_unflattened[1][3] = a[255:224];
  assign a_unflattened[2][0] = a[287:256];
  assign a_unflattened[2][1] = a[319:288];
  assign a_unflattened[2][2] = a[351:320];
  assign a_unflattened[2][3] = a[383:352];
  assign a_unflattened[3][0] = a[415:384];
  assign a_unflattened[3][1] = a[447:416];
  assign a_unflattened[3][2] = a[479:448];
  assign a_unflattened[3][3] = a[511:480];
  wire [31:0] b_unflattened[4][4];
  assign b_unflattened[0][0] = b[31:0];
  assign b_unflattened[0][1] = b[63:32];
  assign b_unflattened[0][2] = b[95:64];
  assign b_unflattened[0][3] = b[127:96];
  assign b_unflattened[1][0] = b[159:128];
  assign b_unflattened[1][1] = b[191:160];
  assign b_unflattened[1][2] = b[223:192];
  assign b_unflattened[1][3] = b[255:224];
  assign b_unflattened[2][0] = b[287:256];
  assign b_unflattened[2][1] = b[319:288];
  assign b_unflattened[2][2] = b[351:320];
  assign b_unflattened[2][3] = b[383:352];
  assign b_unflattened[3][0] = b[415:384];
  assign b_unflattened[3][1] = b[447:416];
  assign b_unflattened[3][2] = b[479:448];
  assign b_unflattened[3][3] = b[511:480];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [31:0] p0_a[4][4];
  reg [31:0] p0_b[4][4];
  always_ff @ (posedge clk) begin
    p0_a <= a_unflattened;
    p0_b <= b_unflattened;
  end

  // ===== Pipe stage 1:
  wire [31:0] p1_array_index_663_comb;
  wire [31:0] p1_array_index_664_comb;
  wire [31:0] p1_array_index_665_comb;
  wire [31:0] p1_array_index_666_comb;
  wire [31:0] p1_array_index_667_comb;
  wire [31:0] p1_array_index_668_comb;
  wire [31:0] p1_array_index_669_comb;
  wire [31:0] p1_array_index_670_comb;
  wire [31:0] p1_array_index_671_comb;
  wire [31:0] p1_array_index_672_comb;
  wire [31:0] p1_array_index_673_comb;
  wire [31:0] p1_array_index_674_comb;
  wire [31:0] p1_array_index_675_comb;
  wire [31:0] p1_array_index_676_comb;
  wire [31:0] p1_array_index_677_comb;
  wire [31:0] p1_array_index_678_comb;
  wire [31:0] p1_array_index_679_comb;
  wire [31:0] p1_array_index_680_comb;
  wire [31:0] p1_array_index_681_comb;
  wire [31:0] p1_array_index_682_comb;
  wire [31:0] p1_array_index_683_comb;
  wire [31:0] p1_array_index_684_comb;
  wire [31:0] p1_array_index_685_comb;
  wire [31:0] p1_array_index_686_comb;
  wire [31:0] p1_array_index_687_comb;
  wire [31:0] p1_array_index_688_comb;
  wire [31:0] p1_array_index_689_comb;
  wire [31:0] p1_array_index_690_comb;
  wire [31:0] p1_array_index_691_comb;
  wire [31:0] p1_array_index_692_comb;
  wire [31:0] p1_array_index_693_comb;
  wire [31:0] p1_array_index_694_comb;
  wire [31:0] p1_smul_695_comb;
  wire [31:0] p1_smul_696_comb;
  wire [31:0] p1_smul_697_comb;
  wire [31:0] p1_smul_698_comb;
  wire [31:0] p1_smul_699_comb;
  wire [31:0] p1_smul_700_comb;
  wire [31:0] p1_smul_701_comb;
  wire [31:0] p1_smul_702_comb;
  wire [31:0] p1_smul_703_comb;
  wire [31:0] p1_smul_704_comb;
  wire [31:0] p1_smul_705_comb;
  wire [31:0] p1_smul_706_comb;
  wire [31:0] p1_smul_707_comb;
  wire [31:0] p1_smul_708_comb;
  wire [31:0] p1_smul_709_comb;
  wire [31:0] p1_smul_710_comb;
  wire [31:0] p1_smul_711_comb;
  wire [31:0] p1_smul_712_comb;
  wire [31:0] p1_smul_713_comb;
  wire [31:0] p1_smul_714_comb;
  wire [31:0] p1_smul_715_comb;
  wire [31:0] p1_smul_716_comb;
  wire [31:0] p1_smul_717_comb;
  wire [31:0] p1_smul_718_comb;
  wire [31:0] p1_smul_719_comb;
  wire [31:0] p1_smul_720_comb;
  wire [31:0] p1_smul_721_comb;
  wire [31:0] p1_smul_722_comb;
  wire [31:0] p1_smul_723_comb;
  wire [31:0] p1_smul_724_comb;
  wire [31:0] p1_smul_725_comb;
  wire [31:0] p1_smul_726_comb;
  wire [31:0] p1_smul_727_comb;
  wire [31:0] p1_smul_728_comb;
  wire [31:0] p1_smul_729_comb;
  wire [31:0] p1_smul_730_comb;
  wire [31:0] p1_smul_731_comb;
  wire [31:0] p1_smul_732_comb;
  wire [31:0] p1_smul_733_comb;
  wire [31:0] p1_smul_734_comb;
  wire [31:0] p1_smul_735_comb;
  wire [31:0] p1_smul_736_comb;
  wire [31:0] p1_smul_737_comb;
  wire [31:0] p1_smul_738_comb;
  wire [31:0] p1_smul_739_comb;
  wire [31:0] p1_smul_740_comb;
  wire [31:0] p1_smul_741_comb;
  wire [31:0] p1_smul_742_comb;
  wire [31:0] p1_smul_743_comb;
  wire [31:0] p1_smul_744_comb;
  wire [31:0] p1_smul_745_comb;
  wire [31:0] p1_smul_746_comb;
  wire [31:0] p1_smul_747_comb;
  wire [31:0] p1_smul_748_comb;
  wire [31:0] p1_smul_749_comb;
  wire [31:0] p1_smul_750_comb;
  wire [31:0] p1_smul_751_comb;
  wire [31:0] p1_smul_752_comb;
  wire [31:0] p1_smul_753_comb;
  wire [31:0] p1_smul_754_comb;
  wire [31:0] p1_smul_755_comb;
  wire [31:0] p1_smul_756_comb;
  wire [31:0] p1_smul_757_comb;
  wire [31:0] p1_smul_758_comb;
  wire [31:0] p1_dot_associative_element_comb;
  wire [31:0] p1_dot_associative_element__1_comb;
  wire [31:0] p1_dot_associative_element__2_comb;
  wire [31:0] p1_dot_associative_element__3_comb;
  wire [31:0] p1_dot_associative_element__4_comb;
  wire [31:0] p1_dot_associative_element__5_comb;
  wire [31:0] p1_dot_associative_element__6_comb;
  wire [31:0] p1_dot_associative_element__7_comb;
  wire [31:0] p1_dot_associative_element__8_comb;
  wire [31:0] p1_dot_associative_element__9_comb;
  wire [31:0] p1_dot_associative_element__10_comb;
  wire [31:0] p1_dot_associative_element__11_comb;
  wire [31:0] p1_dot_associative_element__12_comb;
  wire [31:0] p1_dot_associative_element__13_comb;
  wire [31:0] p1_dot_associative_element__14_comb;
  wire [31:0] p1_dot_associative_element__15_comb;
  wire [31:0] p1_dot_associative_element__16_comb;
  wire [31:0] p1_dot_associative_element__17_comb;
  wire [31:0] p1_dot_associative_element__18_comb;
  wire [31:0] p1_dot_associative_element__19_comb;
  wire [31:0] p1_dot_associative_element__20_comb;
  wire [31:0] p1_dot_associative_element__21_comb;
  wire [31:0] p1_dot_associative_element__22_comb;
  wire [31:0] p1_dot_associative_element__23_comb;
  wire [31:0] p1_dot_associative_element__24_comb;
  wire [31:0] p1_dot_associative_element__25_comb;
  wire [31:0] p1_dot_associative_element__26_comb;
  wire [31:0] p1_dot_associative_element__27_comb;
  wire [31:0] p1_dot_associative_element__28_comb;
  wire [31:0] p1_dot_associative_element__29_comb;
  wire [31:0] p1_dot_associative_element__30_comb;
  wire [31:0] p1_dot_associative_element__31_comb;
  wire [31:0] p1_dot_comb;
  wire [31:0] p1_dot__1_comb;
  wire [31:0] p1_dot__2_comb;
  wire [31:0] p1_dot__3_comb;
  wire [31:0] p1_dot__4_comb;
  wire [31:0] p1_dot__5_comb;
  wire [31:0] p1_dot__6_comb;
  wire [31:0] p1_dot__7_comb;
  wire [31:0] p1_dot__8_comb;
  wire [31:0] p1_dot__9_comb;
  wire [31:0] p1_dot__10_comb;
  wire [31:0] p1_dot__11_comb;
  wire [31:0] p1_dot__12_comb;
  wire [31:0] p1_dot__13_comb;
  wire [31:0] p1_dot__14_comb;
  wire [31:0] p1_dot__15_comb;
  wire [31:0] p1_row_comb[4];
  wire [31:0] p1_row__1_comb[4];
  wire [31:0] p1_row__2_comb[4];
  wire [31:0] p1_row__3_comb[4];
  wire [31:0] p1_array_811_comb[4][4];
  assign p1_array_index_663_comb = p0_a[2'h0][2'h0];
  assign p1_array_index_664_comb = p0_b[2'h0][2'h0];
  assign p1_array_index_665_comb = p0_a[2'h0][2'h1];
  assign p1_array_index_666_comb = p0_b[2'h1][2'h0];
  assign p1_array_index_667_comb = p0_a[2'h0][2'h2];
  assign p1_array_index_668_comb = p0_b[2'h2][2'h0];
  assign p1_array_index_669_comb = p0_a[2'h0][2'h3];
  assign p1_array_index_670_comb = p0_b[2'h3][2'h0];
  assign p1_array_index_671_comb = p0_b[2'h0][2'h1];
  assign p1_array_index_672_comb = p0_b[2'h1][2'h1];
  assign p1_array_index_673_comb = p0_b[2'h2][2'h1];
  assign p1_array_index_674_comb = p0_b[2'h3][2'h1];
  assign p1_array_index_675_comb = p0_b[2'h0][2'h2];
  assign p1_array_index_676_comb = p0_b[2'h1][2'h2];
  assign p1_array_index_677_comb = p0_b[2'h2][2'h2];
  assign p1_array_index_678_comb = p0_b[2'h3][2'h2];
  assign p1_array_index_679_comb = p0_b[2'h0][2'h3];
  assign p1_array_index_680_comb = p0_b[2'h1][2'h3];
  assign p1_array_index_681_comb = p0_b[2'h2][2'h3];
  assign p1_array_index_682_comb = p0_b[2'h3][2'h3];
  assign p1_array_index_683_comb = p0_a[2'h1][2'h0];
  assign p1_array_index_684_comb = p0_a[2'h1][2'h1];
  assign p1_array_index_685_comb = p0_a[2'h1][2'h2];
  assign p1_array_index_686_comb = p0_a[2'h1][2'h3];
  assign p1_array_index_687_comb = p0_a[2'h2][2'h0];
  assign p1_array_index_688_comb = p0_a[2'h2][2'h1];
  assign p1_array_index_689_comb = p0_a[2'h2][2'h2];
  assign p1_array_index_690_comb = p0_a[2'h2][2'h3];
  assign p1_array_index_691_comb = p0_a[2'h3][2'h0];
  assign p1_array_index_692_comb = p0_a[2'h3][2'h1];
  assign p1_array_index_693_comb = p0_a[2'h3][2'h2];
  assign p1_array_index_694_comb = p0_a[2'h3][2'h3];
  assign p1_smul_695_comb = smul32b_32b_x_32b(p1_array_index_663_comb, p1_array_index_664_comb);
  assign p1_smul_696_comb = smul32b_32b_x_32b(p1_array_index_665_comb, p1_array_index_666_comb);
  assign p1_smul_697_comb = smul32b_32b_x_32b(p1_array_index_667_comb, p1_array_index_668_comb);
  assign p1_smul_698_comb = smul32b_32b_x_32b(p1_array_index_669_comb, p1_array_index_670_comb);
  assign p1_smul_699_comb = smul32b_32b_x_32b(p1_array_index_663_comb, p1_array_index_671_comb);
  assign p1_smul_700_comb = smul32b_32b_x_32b(p1_array_index_665_comb, p1_array_index_672_comb);
  assign p1_smul_701_comb = smul32b_32b_x_32b(p1_array_index_667_comb, p1_array_index_673_comb);
  assign p1_smul_702_comb = smul32b_32b_x_32b(p1_array_index_669_comb, p1_array_index_674_comb);
  assign p1_smul_703_comb = smul32b_32b_x_32b(p1_array_index_663_comb, p1_array_index_675_comb);
  assign p1_smul_704_comb = smul32b_32b_x_32b(p1_array_index_665_comb, p1_array_index_676_comb);
  assign p1_smul_705_comb = smul32b_32b_x_32b(p1_array_index_667_comb, p1_array_index_677_comb);
  assign p1_smul_706_comb = smul32b_32b_x_32b(p1_array_index_669_comb, p1_array_index_678_comb);
  assign p1_smul_707_comb = smul32b_32b_x_32b(p1_array_index_663_comb, p1_array_index_679_comb);
  assign p1_smul_708_comb = smul32b_32b_x_32b(p1_array_index_665_comb, p1_array_index_680_comb);
  assign p1_smul_709_comb = smul32b_32b_x_32b(p1_array_index_667_comb, p1_array_index_681_comb);
  assign p1_smul_710_comb = smul32b_32b_x_32b(p1_array_index_669_comb, p1_array_index_682_comb);
  assign p1_smul_711_comb = smul32b_32b_x_32b(p1_array_index_683_comb, p1_array_index_664_comb);
  assign p1_smul_712_comb = smul32b_32b_x_32b(p1_array_index_684_comb, p1_array_index_666_comb);
  assign p1_smul_713_comb = smul32b_32b_x_32b(p1_array_index_685_comb, p1_array_index_668_comb);
  assign p1_smul_714_comb = smul32b_32b_x_32b(p1_array_index_686_comb, p1_array_index_670_comb);
  assign p1_smul_715_comb = smul32b_32b_x_32b(p1_array_index_683_comb, p1_array_index_671_comb);
  assign p1_smul_716_comb = smul32b_32b_x_32b(p1_array_index_684_comb, p1_array_index_672_comb);
  assign p1_smul_717_comb = smul32b_32b_x_32b(p1_array_index_685_comb, p1_array_index_673_comb);
  assign p1_smul_718_comb = smul32b_32b_x_32b(p1_array_index_686_comb, p1_array_index_674_comb);
  assign p1_smul_719_comb = smul32b_32b_x_32b(p1_array_index_683_comb, p1_array_index_675_comb);
  assign p1_smul_720_comb = smul32b_32b_x_32b(p1_array_index_684_comb, p1_array_index_676_comb);
  assign p1_smul_721_comb = smul32b_32b_x_32b(p1_array_index_685_comb, p1_array_index_677_comb);
  assign p1_smul_722_comb = smul32b_32b_x_32b(p1_array_index_686_comb, p1_array_index_678_comb);
  assign p1_smul_723_comb = smul32b_32b_x_32b(p1_array_index_683_comb, p1_array_index_679_comb);
  assign p1_smul_724_comb = smul32b_32b_x_32b(p1_array_index_684_comb, p1_array_index_680_comb);
  assign p1_smul_725_comb = smul32b_32b_x_32b(p1_array_index_685_comb, p1_array_index_681_comb);
  assign p1_smul_726_comb = smul32b_32b_x_32b(p1_array_index_686_comb, p1_array_index_682_comb);
  assign p1_smul_727_comb = smul32b_32b_x_32b(p1_array_index_687_comb, p1_array_index_664_comb);
  assign p1_smul_728_comb = smul32b_32b_x_32b(p1_array_index_688_comb, p1_array_index_666_comb);
  assign p1_smul_729_comb = smul32b_32b_x_32b(p1_array_index_689_comb, p1_array_index_668_comb);
  assign p1_smul_730_comb = smul32b_32b_x_32b(p1_array_index_690_comb, p1_array_index_670_comb);
  assign p1_smul_731_comb = smul32b_32b_x_32b(p1_array_index_687_comb, p1_array_index_671_comb);
  assign p1_smul_732_comb = smul32b_32b_x_32b(p1_array_index_688_comb, p1_array_index_672_comb);
  assign p1_smul_733_comb = smul32b_32b_x_32b(p1_array_index_689_comb, p1_array_index_673_comb);
  assign p1_smul_734_comb = smul32b_32b_x_32b(p1_array_index_690_comb, p1_array_index_674_comb);
  assign p1_smul_735_comb = smul32b_32b_x_32b(p1_array_index_687_comb, p1_array_index_675_comb);
  assign p1_smul_736_comb = smul32b_32b_x_32b(p1_array_index_688_comb, p1_array_index_676_comb);
  assign p1_smul_737_comb = smul32b_32b_x_32b(p1_array_index_689_comb, p1_array_index_677_comb);
  assign p1_smul_738_comb = smul32b_32b_x_32b(p1_array_index_690_comb, p1_array_index_678_comb);
  assign p1_smul_739_comb = smul32b_32b_x_32b(p1_array_index_687_comb, p1_array_index_679_comb);
  assign p1_smul_740_comb = smul32b_32b_x_32b(p1_array_index_688_comb, p1_array_index_680_comb);
  assign p1_smul_741_comb = smul32b_32b_x_32b(p1_array_index_689_comb, p1_array_index_681_comb);
  assign p1_smul_742_comb = smul32b_32b_x_32b(p1_array_index_690_comb, p1_array_index_682_comb);
  assign p1_smul_743_comb = smul32b_32b_x_32b(p1_array_index_691_comb, p1_array_index_664_comb);
  assign p1_smul_744_comb = smul32b_32b_x_32b(p1_array_index_692_comb, p1_array_index_666_comb);
  assign p1_smul_745_comb = smul32b_32b_x_32b(p1_array_index_693_comb, p1_array_index_668_comb);
  assign p1_smul_746_comb = smul32b_32b_x_32b(p1_array_index_694_comb, p1_array_index_670_comb);
  assign p1_smul_747_comb = smul32b_32b_x_32b(p1_array_index_691_comb, p1_array_index_671_comb);
  assign p1_smul_748_comb = smul32b_32b_x_32b(p1_array_index_692_comb, p1_array_index_672_comb);
  assign p1_smul_749_comb = smul32b_32b_x_32b(p1_array_index_693_comb, p1_array_index_673_comb);
  assign p1_smul_750_comb = smul32b_32b_x_32b(p1_array_index_694_comb, p1_array_index_674_comb);
  assign p1_smul_751_comb = smul32b_32b_x_32b(p1_array_index_691_comb, p1_array_index_675_comb);
  assign p1_smul_752_comb = smul32b_32b_x_32b(p1_array_index_692_comb, p1_array_index_676_comb);
  assign p1_smul_753_comb = smul32b_32b_x_32b(p1_array_index_693_comb, p1_array_index_677_comb);
  assign p1_smul_754_comb = smul32b_32b_x_32b(p1_array_index_694_comb, p1_array_index_678_comb);
  assign p1_smul_755_comb = smul32b_32b_x_32b(p1_array_index_691_comb, p1_array_index_679_comb);
  assign p1_smul_756_comb = smul32b_32b_x_32b(p1_array_index_692_comb, p1_array_index_680_comb);
  assign p1_smul_757_comb = smul32b_32b_x_32b(p1_array_index_693_comb, p1_array_index_681_comb);
  assign p1_smul_758_comb = smul32b_32b_x_32b(p1_array_index_694_comb, p1_array_index_682_comb);
  assign p1_dot_associative_element_comb = p1_smul_695_comb + p1_smul_696_comb;
  assign p1_dot_associative_element__1_comb = p1_smul_697_comb + p1_smul_698_comb;
  assign p1_dot_associative_element__2_comb = p1_smul_699_comb + p1_smul_700_comb;
  assign p1_dot_associative_element__3_comb = p1_smul_701_comb + p1_smul_702_comb;
  assign p1_dot_associative_element__4_comb = p1_smul_703_comb + p1_smul_704_comb;
  assign p1_dot_associative_element__5_comb = p1_smul_705_comb + p1_smul_706_comb;
  assign p1_dot_associative_element__6_comb = p1_smul_707_comb + p1_smul_708_comb;
  assign p1_dot_associative_element__7_comb = p1_smul_709_comb + p1_smul_710_comb;
  assign p1_dot_associative_element__8_comb = p1_smul_711_comb + p1_smul_712_comb;
  assign p1_dot_associative_element__9_comb = p1_smul_713_comb + p1_smul_714_comb;
  assign p1_dot_associative_element__10_comb = p1_smul_715_comb + p1_smul_716_comb;
  assign p1_dot_associative_element__11_comb = p1_smul_717_comb + p1_smul_718_comb;
  assign p1_dot_associative_element__12_comb = p1_smul_719_comb + p1_smul_720_comb;
  assign p1_dot_associative_element__13_comb = p1_smul_721_comb + p1_smul_722_comb;
  assign p1_dot_associative_element__14_comb = p1_smul_723_comb + p1_smul_724_comb;
  assign p1_dot_associative_element__15_comb = p1_smul_725_comb + p1_smul_726_comb;
  assign p1_dot_associative_element__16_comb = p1_smul_727_comb + p1_smul_728_comb;
  assign p1_dot_associative_element__17_comb = p1_smul_729_comb + p1_smul_730_comb;
  assign p1_dot_associative_element__18_comb = p1_smul_731_comb + p1_smul_732_comb;
  assign p1_dot_associative_element__19_comb = p1_smul_733_comb + p1_smul_734_comb;
  assign p1_dot_associative_element__20_comb = p1_smul_735_comb + p1_smul_736_comb;
  assign p1_dot_associative_element__21_comb = p1_smul_737_comb + p1_smul_738_comb;
  assign p1_dot_associative_element__22_comb = p1_smul_739_comb + p1_smul_740_comb;
  assign p1_dot_associative_element__23_comb = p1_smul_741_comb + p1_smul_742_comb;
  assign p1_dot_associative_element__24_comb = p1_smul_743_comb + p1_smul_744_comb;
  assign p1_dot_associative_element__25_comb = p1_smul_745_comb + p1_smul_746_comb;
  assign p1_dot_associative_element__26_comb = p1_smul_747_comb + p1_smul_748_comb;
  assign p1_dot_associative_element__27_comb = p1_smul_749_comb + p1_smul_750_comb;
  assign p1_dot_associative_element__28_comb = p1_smul_751_comb + p1_smul_752_comb;
  assign p1_dot_associative_element__29_comb = p1_smul_753_comb + p1_smul_754_comb;
  assign p1_dot_associative_element__30_comb = p1_smul_755_comb + p1_smul_756_comb;
  assign p1_dot_associative_element__31_comb = p1_smul_757_comb + p1_smul_758_comb;
  assign p1_dot_comb = p1_dot_associative_element_comb + p1_dot_associative_element__1_comb;
  assign p1_dot__1_comb = p1_dot_associative_element__2_comb + p1_dot_associative_element__3_comb;
  assign p1_dot__2_comb = p1_dot_associative_element__4_comb + p1_dot_associative_element__5_comb;
  assign p1_dot__3_comb = p1_dot_associative_element__6_comb + p1_dot_associative_element__7_comb;
  assign p1_dot__4_comb = p1_dot_associative_element__8_comb + p1_dot_associative_element__9_comb;
  assign p1_dot__5_comb = p1_dot_associative_element__10_comb + p1_dot_associative_element__11_comb;
  assign p1_dot__6_comb = p1_dot_associative_element__12_comb + p1_dot_associative_element__13_comb;
  assign p1_dot__7_comb = p1_dot_associative_element__14_comb + p1_dot_associative_element__15_comb;
  assign p1_dot__8_comb = p1_dot_associative_element__16_comb + p1_dot_associative_element__17_comb;
  assign p1_dot__9_comb = p1_dot_associative_element__18_comb + p1_dot_associative_element__19_comb;
  assign p1_dot__10_comb = p1_dot_associative_element__20_comb + p1_dot_associative_element__21_comb;
  assign p1_dot__11_comb = p1_dot_associative_element__22_comb + p1_dot_associative_element__23_comb;
  assign p1_dot__12_comb = p1_dot_associative_element__24_comb + p1_dot_associative_element__25_comb;
  assign p1_dot__13_comb = p1_dot_associative_element__26_comb + p1_dot_associative_element__27_comb;
  assign p1_dot__14_comb = p1_dot_associative_element__28_comb + p1_dot_associative_element__29_comb;
  assign p1_dot__15_comb = p1_dot_associative_element__30_comb + p1_dot_associative_element__31_comb;
  assign p1_row_comb[0] = p1_dot_comb;
  assign p1_row_comb[1] = p1_dot__1_comb;
  assign p1_row_comb[2] = p1_dot__2_comb;
  assign p1_row_comb[3] = p1_dot__3_comb;
  assign p1_row__1_comb[0] = p1_dot__4_comb;
  assign p1_row__1_comb[1] = p1_dot__5_comb;
  assign p1_row__1_comb[2] = p1_dot__6_comb;
  assign p1_row__1_comb[3] = p1_dot__7_comb;
  assign p1_row__2_comb[0] = p1_dot__8_comb;
  assign p1_row__2_comb[1] = p1_dot__9_comb;
  assign p1_row__2_comb[2] = p1_dot__10_comb;
  assign p1_row__2_comb[3] = p1_dot__11_comb;
  assign p1_row__3_comb[0] = p1_dot__12_comb;
  assign p1_row__3_comb[1] = p1_dot__13_comb;
  assign p1_row__3_comb[2] = p1_dot__14_comb;
  assign p1_row__3_comb[3] = p1_dot__15_comb;
  assign p1_array_811_comb[0] = p1_row_comb;
  assign p1_array_811_comb[1] = p1_row__1_comb;
  assign p1_array_811_comb[2] = p1_row__2_comb;
  assign p1_array_811_comb[3] = p1_row__3_comb;

  // Registers for pipe stage 1:
  reg [31:0] p1_array_811[4][4];
  always_ff @ (posedge clk) begin
    p1_array_811 <= p1_array_811_comb;
  end
  assign out = {{p1_array_811[3][3], p1_array_811[3][2], p1_array_811[3][1], p1_array_811[3][0]}, {p1_array_811[2][3], p1_array_811[2][2], p1_array_811[2][1], p1_array_811[2][0]}, {p1_array_811[1][3], p1_array_811[1][2], p1_array_811[1][1], p1_array_811[1][0]}, {p1_array_811[0][3], p1_array_811[0][2], p1_array_811[0][1], p1_array_811[0][0]}};
endmodule
