module __mm__mm_0_next(
  input wire clk,
  input wire rst,
  input wire mm__done_rdy,
  input wire mm__go,
  input wire mm__go_vld,
  input wire mm__mem0__read_req_rdy,
  input wire [31:0] mm__mem0__read_resp,
  input wire mm__mem0__read_resp_vld,
  input wire mm__mem1__read_req_rdy,
  input wire [31:0] mm__mem1__read_resp,
  input wire mm__mem1__read_resp_vld,
  input wire mm__mem2__write_req_rdy,
  input wire mm__mem2__write_resp_vld,
  output wire mm__done,
  output wire mm__done_vld,
  output wire mm__go_rdy,
  output wire [3:0] mm__mem0__read_req,
  output wire mm__mem0__read_req_vld,
  output wire mm__mem0__read_resp_rdy,
  output wire [3:0] mm__mem1__read_req,
  output wire mm__mem1__read_req_vld,
  output wire mm__mem1__read_resp_rdy,
  output wire [35:0] mm__mem2__write_req,
  output wire mm__mem2__write_req_vld,
  output wire mm__mem2__write_resp_rdy
);
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [31:0] smul32b_32b_x_32b (input reg [31:0] lhs, input reg [31:0] rhs);
    reg signed [31:0] signed_lhs;
    reg signed [31:0] signed_rhs;
    reg signed [31:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul32b_32b_x_32b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  wire [31:0] __mm__mem0__read_resp_reg_init = 32'h0000_0000;
  wire [31:0] __mm__mem1__read_resp_reg_init = 32'h0000_0000;
  wire [3:0] __mm__mem0__read_req_reg_init = 4'h0;
  wire [3:0] __mm__mem1__read_req_reg_init = 4'h0;
  wire [35:0] __mm__mem2__write_req_reg_init = {4'h0, 32'h0000_0000};
  reg [31:0] ____state_2;
  reg [31:0] ____state_1;
  reg [1:0] ____state_3;
  reg ____state_4;
  reg p0_or_679;
  reg p0_slt_687;
  reg [3:0] p0_tmp21;
  reg p0_and_712;
  reg p0_tmp27;
  reg p0_and_701;
  reg p0_and_702;
  reg p1_or_679;
  reg p1_slt_687;
  reg [3:0] p1_tmp21;
  reg p1_and_712;
  reg p1_tmp27;
  reg p1_and_701;
  reg p1_and_702;
  reg p2_or_679;
  reg p2_slt_687;
  reg [3:0] p2_tmp21;
  reg p2_and_712;
  reg p2_tmp27;
  reg p2_and_701;
  reg p2_and_702;
  reg p3_or_679;
  reg p3_slt_687;
  reg [3:0] p3_tmp21;
  reg p3_and_712;
  reg p3_tmp27;
  reg p3_and_701;
  reg p3_and_702;
  reg [31:0] ____state_0;
  reg p4_and_712;
  reg p4_tmp27;
  reg p5_and_712;
  reg p5_tmp27;
  reg p6_and_712;
  reg p6_tmp27;
  reg p7_and_712;
  reg p7_tmp27;
  reg p0_valid;
  reg p1_valid;
  reg p2_valid;
  reg p3_valid;
  reg p4_valid;
  reg p5_valid;
  reg p6_valid;
  reg p7_valid;
  reg __mm__mem0__read_req_has_been_sent_reg;
  reg __mm__mem1__read_req_has_been_sent_reg;
  reg __mm__mem2__write_req_has_been_sent_reg;
  reg __mm__done_has_been_sent_reg;
  reg __mm__go_reg;
  reg __mm__go_valid_reg;
  reg [31:0] __mm__mem0__read_resp_reg;
  reg __mm__mem0__read_resp_valid_reg;
  reg [31:0] __mm__mem1__read_resp_reg;
  reg __mm__mem1__read_resp_valid_reg;
  reg __mm__mem2__write_resp_valid_reg;
  reg [3:0] __mm__mem0__read_req_reg;
  reg __mm__mem0__read_req_valid_reg;
  reg [3:0] __mm__mem1__read_req_reg;
  reg __mm__mem1__read_req_valid_reg;
  reg [35:0] __mm__mem2__write_req_reg;
  reg __mm__mem2__write_req_valid_reg;
  reg __mm__done_reg;
  reg __mm__done_valid_reg;
  wire or_895;
  wire __mm__done_vld_buf;
  wire __mm__done_not_has_been_sent;
  wire mm__done_valid_inv;
  wire __mm__done_valid_and_not_has_been_sent;
  wire mm__done_valid_load_en;
  wire mm__done_load_en;
  wire or_1229;
  wire p8_stage_done;
  wire p8_not_valid;
  wire p7_enable;
  wire p7_data_enable;
  wire p7_not_valid;
  wire p6_enable;
  wire p6_data_enable;
  wire p6_not_valid;
  wire p5_enable;
  wire p5_data_enable;
  wire p5_not_valid;
  wire p4_all_active_inputs_valid;
  wire p4_enable;
  wire __mm__mem2__write_req_vld_buf;
  wire __mm__mem2__write_req_not_has_been_sent;
  wire mm__mem2__write_req_valid_inv;
  wire __mm__mem2__write_req_valid_and_not_has_been_sent;
  wire mm__mem2__write_req_valid_load_en;
  wire mm__mem2__write_req_load_en;
  wire or_1228;
  wire p4_stage_done;
  wire p4_data_enable;
  wire p4_not_valid;
  wire p3_enable;
  wire p3_data_enable;
  wire p3_not_valid;
  wire p2_enable;
  wire p2_data_enable;
  wire p2_not_valid;
  wire p1_enable;
  wire p1_data_enable;
  wire p1_not_valid;
  wire or_886;
  wire p0_enable;
  wire __mm__mem0__read_req_vld_buf;
  wire __mm__mem0__read_req_not_has_been_sent;
  wire mm__mem0__read_req_valid_inv;
  wire __mm__mem1__read_req_not_has_been_sent;
  wire mm__mem1__read_req_valid_inv;
  wire [2:0] add_680;
  wire [31:0] add_681;
  wire [31:0] add_682;
  wire __mm__mem0__read_req_valid_and_not_has_been_sent;
  wire mm__mem0__read_req_valid_load_en;
  wire __mm__mem1__read_req_valid_and_not_has_been_sent;
  wire mm__mem1__read_req_valid_load_en;
  wire tmp20;
  wire sge_685;
  wire sge_686;
  wire slt_687;
  wire slt_688;
  wire mm__mem0__read_req_load_en;
  wire mm__mem1__read_req_load_en;
  wire nand_690;
  wire __mm__mem0__read_req_has_sent_or_is_ready;
  wire __mm__mem1__read_req_has_sent_or_is_ready;
  wire tmp27;
  wire and_701;
  wire and_702;
  wire nor_703;
  wire tmp25;
  wire nor_705;
  wire p0_all_active_outputs_ready;
  wire [2:0] ____state_0__next_value_predicates;
  wire [1:0] ____state_1__next_value_predicates;
  wire [1:0] ____state_2__next_value_predicates;
  wire [1:0] ____state_3__next_value_predicates;
  wire p0_stage_done;
  wire [3:0] one_hot_714;
  wire [2:0] one_hot_715;
  wire [2:0] one_hot_716;
  wire [2:0] one_hot_717;
  wire [31:0] tmp6_data;
  wire [31:0] tmp10_data;
  wire p0_data_enable;
  wire mm__go_select;
  wire [31:0] tmp3;
  wire [31:0] tmp15;
  wire mm__go_valid_inv;
  wire mm__mem0__read_resp_valid_inv;
  wire mm__mem1__read_resp_valid_inv;
  wire mm__mem2__write_resp_valid_inv;
  wire [1:0] tmp4__2;
  wire and_1035;
  wire and_1036;
  wire and_1037;
  wire and_1043;
  wire and_1044;
  wire and_1050;
  wire and_1051;
  wire and_1058;
  wire and_1059;
  wire [1:0] add_667;
  wire [31:0] tmp17;
  wire mm__go_valid_load_en;
  wire mm__mem0__read_resp_valid_load_en;
  wire mm__mem1__read_resp_valid_load_en;
  wire mm__mem2__write_resp_valid_load_en;
  wire ____state_0__at_most_one_next_value;
  wire ____state_1__at_most_one_next_value;
  wire ____state_2__at_most_one_next_value;
  wire ____state_3__at_most_one_next_value;
  wire [1:0] add_699;
  wire [2:0] concat_1039;
  wire [31:0] tmp2;
  wire [1:0] concat_1046;
  wire [1:0] concat_1053;
  wire tmp1;
  wire [1:0] concat_1060;
  wire [1:0] unexpand_for_next_value_158_3_case_1;
  wire [1:0] unexpand_for_next_value_158_3_case_0;
  wire __mm__mem0__read_req_valid_and_all_active_outputs_ready;
  wire __mm__mem0__read_req_valid_and_ready_txfr;
  wire __mm__mem1__read_req_valid_and_ready_txfr;
  wire __mm__mem2__write_req_valid_and_all_active_outputs_ready;
  wire __mm__mem2__write_req_valid_and_ready_txfr;
  wire __mm__done_valid_and_all_active_outputs_ready;
  wire __mm__done_valid_and_ready_txfr;
  wire [3:0] tmp4;
  wire [3:0] tmp8;
  wire [31:0] tmp18;
  wire mm__go_load_en;
  wire mm__mem0__read_resp_load_en;
  wire mm__mem1__read_resp_load_en;
  wire mm__mem2__write_resp_load_en;
  wire or_1221;
  wire or_1223;
  wire or_1225;
  wire or_1227;
  wire or_679;
  wire [3:0] tmp21;
  wire and_712;
  wire [31:0] one_hot_sel_1040;
  wire or_1041;
  wire [31:0] one_hot_sel_1047;
  wire or_1048;
  wire [31:0] one_hot_sel_1054;
  wire or_1055;
  wire tmp32;
  wire [1:0] one_hot_sel_1061;
  wire or_1062;
  wire __mm__mem0__read_req_not_stage_load;
  wire __mm__mem0__read_req_has_been_sent_reg_load_en;
  wire __mm__mem1__read_req_has_been_sent_reg_load_en;
  wire __mm__mem2__write_req_not_stage_load;
  wire __mm__mem2__write_req_has_been_sent_reg_load_en;
  wire __mm__done_not_stage_load;
  wire __mm__done_has_been_sent_reg_load_en;
  wire [3:0] tmp5;
  wire [3:0] tmp9;
  wire [35:0] tmp23;
  wire __mm__done_buf;
  assign or_895 = ~p7_and_712 | __mm__mem2__write_resp_valid_reg;
  assign __mm__done_vld_buf = or_895 & p7_valid & p7_tmp27;
  assign __mm__done_not_has_been_sent = ~__mm__done_has_been_sent_reg;
  assign mm__done_valid_inv = ~__mm__done_valid_reg;
  assign __mm__done_valid_and_not_has_been_sent = __mm__done_vld_buf & __mm__done_not_has_been_sent;
  assign mm__done_valid_load_en = mm__done_rdy | mm__done_valid_inv;
  assign mm__done_load_en = __mm__done_valid_and_not_has_been_sent & mm__done_valid_load_en;
  assign or_1229 = ~p7_tmp27 | mm__done_load_en | __mm__done_has_been_sent_reg;
  assign p8_stage_done = p7_valid & or_895 & or_1229;
  assign p8_not_valid = ~p7_valid;
  assign p7_enable = p8_stage_done | p8_not_valid;
  assign p7_data_enable = p7_enable & p6_valid;
  assign p7_not_valid = ~p6_valid;
  assign p6_enable = p7_data_enable | p7_not_valid;
  assign p6_data_enable = p6_enable & p5_valid;
  assign p6_not_valid = ~p5_valid;
  assign p5_enable = p6_data_enable | p6_not_valid;
  assign p5_data_enable = p5_enable & p4_valid;
  assign p5_not_valid = ~p4_valid;
  assign p4_all_active_inputs_valid = __mm__mem0__read_resp_valid_reg & __mm__mem1__read_resp_valid_reg;
  assign p4_enable = p5_data_enable | p5_not_valid;
  assign __mm__mem2__write_req_vld_buf = p4_all_active_inputs_valid & p3_valid & p4_enable & p3_and_712;
  assign __mm__mem2__write_req_not_has_been_sent = ~__mm__mem2__write_req_has_been_sent_reg;
  assign mm__mem2__write_req_valid_inv = ~__mm__mem2__write_req_valid_reg;
  assign __mm__mem2__write_req_valid_and_not_has_been_sent = __mm__mem2__write_req_vld_buf & __mm__mem2__write_req_not_has_been_sent;
  assign mm__mem2__write_req_valid_load_en = mm__mem2__write_req_rdy | mm__mem2__write_req_valid_inv;
  assign mm__mem2__write_req_load_en = __mm__mem2__write_req_valid_and_not_has_been_sent & mm__mem2__write_req_valid_load_en;
  assign or_1228 = ~p3_and_712 | mm__mem2__write_req_load_en | __mm__mem2__write_req_has_been_sent_reg;
  assign p4_stage_done = p3_valid & p4_all_active_inputs_valid & or_1228;
  assign p4_data_enable = p4_enable & p4_stage_done;
  assign p4_not_valid = ~p3_valid;
  assign p3_enable = p4_data_enable | p4_not_valid;
  assign p3_data_enable = p3_enable & p2_valid;
  assign p3_not_valid = ~p2_valid;
  assign p2_enable = p3_data_enable | p3_not_valid;
  assign p2_data_enable = p2_enable & p1_valid;
  assign p2_not_valid = ~p1_valid;
  assign p1_enable = p2_data_enable | p2_not_valid;
  assign p1_data_enable = p1_enable & p0_valid;
  assign p1_not_valid = ~p0_valid;
  assign or_886 = ____state_4 | __mm__go_valid_reg;
  assign p0_enable = p1_data_enable | p1_not_valid;
  assign __mm__mem0__read_req_vld_buf = or_886 & p0_enable;
  assign __mm__mem0__read_req_not_has_been_sent = ~__mm__mem0__read_req_has_been_sent_reg;
  assign mm__mem0__read_req_valid_inv = ~__mm__mem0__read_req_valid_reg;
  assign __mm__mem1__read_req_not_has_been_sent = ~__mm__mem1__read_req_has_been_sent_reg;
  assign mm__mem1__read_req_valid_inv = ~__mm__mem1__read_req_valid_reg;
  assign add_680 = {1'h0, ____state_3} + 3'h1;
  assign add_681 = ____state_2 + 32'h0000_0001;
  assign add_682 = ____state_1 + 32'h0000_0001;
  assign __mm__mem0__read_req_valid_and_not_has_been_sent = __mm__mem0__read_req_vld_buf & __mm__mem0__read_req_not_has_been_sent;
  assign mm__mem0__read_req_valid_load_en = mm__mem0__read_req_rdy | mm__mem0__read_req_valid_inv;
  assign __mm__mem1__read_req_valid_and_not_has_been_sent = __mm__mem0__read_req_vld_buf & __mm__mem1__read_req_not_has_been_sent;
  assign mm__mem1__read_req_valid_load_en = mm__mem1__read_req_rdy | mm__mem1__read_req_valid_inv;
  assign tmp20 = add_680[2];
  assign sge_685 = $signed(add_681) >= $signed(32'h0000_0004);
  assign sge_686 = $signed(add_682) >= $signed(32'h0000_0004);
  assign slt_687 = $signed(____state_1) < $signed(32'h0000_0004);
  assign slt_688 = $signed(____state_2) < $signed(32'h0000_0004);
  assign mm__mem0__read_req_load_en = __mm__mem0__read_req_valid_and_not_has_been_sent & mm__mem0__read_req_valid_load_en;
  assign mm__mem1__read_req_load_en = __mm__mem1__read_req_valid_and_not_has_been_sent & mm__mem1__read_req_valid_load_en;
  assign nand_690 = ~(tmp20 & sge_685 & sge_686);
  assign __mm__mem0__read_req_has_sent_or_is_ready = mm__mem0__read_req_load_en | __mm__mem0__read_req_has_been_sent_reg;
  assign __mm__mem1__read_req_has_sent_or_is_ready = mm__mem1__read_req_load_en | __mm__mem1__read_req_has_been_sent_reg;
  assign tmp27 = tmp20 & sge_685 & sge_686;
  assign and_701 = nand_690 & slt_687 & slt_688;
  assign and_702 = nand_690 & ~(slt_687 & slt_688) & slt_688 & ~(____state_3[0] | ____state_3[1]);
  assign nor_703 = ~(~tmp20 | ~sge_685 | sge_686);
  assign tmp25 = tmp20 & sge_685;
  assign nor_705 = ~(~tmp20 | sge_685);
  assign p0_all_active_outputs_ready = __mm__mem0__read_req_has_sent_or_is_ready & __mm__mem1__read_req_has_sent_or_is_ready;
  assign ____state_0__next_value_predicates = {tmp27, and_701, and_702};
  assign ____state_1__next_value_predicates = {tmp27, nor_703};
  assign ____state_2__next_value_predicates = {tmp25, nor_705};
  assign ____state_3__next_value_predicates = {~tmp20, tmp20};
  assign p0_stage_done = or_886 & p0_all_active_outputs_ready;
  assign one_hot_714 = {____state_0__next_value_predicates[2:0] == 3'h0, ____state_0__next_value_predicates[2] && ____state_0__next_value_predicates[1:0] == 2'h0, ____state_0__next_value_predicates[1] && !____state_0__next_value_predicates[0], ____state_0__next_value_predicates[0]};
  assign one_hot_715 = {____state_1__next_value_predicates[1:0] == 2'h0, ____state_1__next_value_predicates[1] && !____state_1__next_value_predicates[0], ____state_1__next_value_predicates[0]};
  assign one_hot_716 = {____state_2__next_value_predicates[1:0] == 2'h0, ____state_2__next_value_predicates[1] && !____state_2__next_value_predicates[0], ____state_2__next_value_predicates[0]};
  assign one_hot_717 = {____state_3__next_value_predicates[1:0] == 2'h0, ____state_3__next_value_predicates[1] && !____state_3__next_value_predicates[0], ____state_3__next_value_predicates[0]};
  assign tmp6_data = __mm__mem0__read_resp_reg[31:0];
  assign tmp10_data = __mm__mem1__read_resp_reg[31:0];
  assign p0_data_enable = p0_enable & p0_stage_done;
  assign mm__go_select = ~____state_4 ? __mm__go_reg : 1'h0;
  assign tmp3 = ____state_0 & {32{p3_or_679}};
  assign tmp15 = smul32b_32b_x_32b(tmp6_data, tmp10_data);
  assign mm__go_valid_inv = ~__mm__go_valid_reg;
  assign mm__mem0__read_resp_valid_inv = ~__mm__mem0__read_resp_valid_reg;
  assign mm__mem1__read_resp_valid_inv = ~__mm__mem1__read_resp_valid_reg;
  assign mm__mem2__write_resp_valid_inv = ~__mm__mem2__write_resp_valid_reg;
  assign tmp4__2 = ____state_1[1:0];
  assign and_1035 = p3_tmp27 & p4_data_enable;
  assign and_1036 = p3_and_701 & p4_data_enable;
  assign and_1037 = p3_and_702 & p4_data_enable;
  assign and_1043 = tmp27 & p0_data_enable;
  assign and_1044 = nor_703 & p0_data_enable;
  assign and_1050 = tmp25 & p0_data_enable;
  assign and_1051 = nor_705 & p0_data_enable;
  assign and_1058 = ~tmp20 & p0_data_enable;
  assign and_1059 = tmp20 & p0_data_enable;
  assign add_667 = ____state_3 + ____state_2[3:2];
  assign tmp17 = tmp3 + tmp15;
  assign mm__go_valid_load_en = p0_data_enable & ~____state_4 | mm__go_valid_inv;
  assign mm__mem0__read_resp_valid_load_en = p4_data_enable | mm__mem0__read_resp_valid_inv;
  assign mm__mem1__read_resp_valid_load_en = p4_data_enable | mm__mem1__read_resp_valid_inv;
  assign mm__mem2__write_resp_valid_load_en = p8_stage_done & p7_and_712 | mm__mem2__write_resp_valid_inv;
  assign ____state_0__at_most_one_next_value = tmp27 == one_hot_714[2] & and_701 == one_hot_714[1] & and_702 == one_hot_714[0];
  assign ____state_1__at_most_one_next_value = tmp27 == one_hot_715[1] & nor_703 == one_hot_715[0];
  assign ____state_2__at_most_one_next_value = tmp25 == one_hot_716[1] & nor_705 == one_hot_716[0];
  assign ____state_3__at_most_one_next_value = ~tmp20 == one_hot_717[1] & tmp20 == one_hot_717[0];
  assign add_699 = tmp4__2 + ____state_2[3:2];
  assign concat_1039 = {and_1035, and_1036, and_1037};
  assign tmp2 = 32'h0000_0000;
  assign concat_1046 = {and_1043, and_1044};
  assign concat_1053 = {and_1050, and_1051};
  assign tmp1 = ~(____state_4 | ~mm__go_select);
  assign concat_1060 = {and_1058, and_1059};
  assign unexpand_for_next_value_158_3_case_1 = 2'h0;
  assign unexpand_for_next_value_158_3_case_0 = add_680[1:0];
  assign __mm__mem0__read_req_valid_and_all_active_outputs_ready = __mm__mem0__read_req_vld_buf & p0_all_active_outputs_ready;
  assign __mm__mem0__read_req_valid_and_ready_txfr = __mm__mem0__read_req_valid_and_not_has_been_sent & mm__mem0__read_req_load_en;
  assign __mm__mem1__read_req_valid_and_ready_txfr = __mm__mem1__read_req_valid_and_not_has_been_sent & mm__mem1__read_req_load_en;
  assign __mm__mem2__write_req_valid_and_all_active_outputs_ready = __mm__mem2__write_req_vld_buf & or_1228;
  assign __mm__mem2__write_req_valid_and_ready_txfr = __mm__mem2__write_req_valid_and_not_has_been_sent & mm__mem2__write_req_load_en;
  assign __mm__done_valid_and_all_active_outputs_ready = __mm__done_vld_buf & or_1229;
  assign __mm__done_valid_and_ready_txfr = __mm__done_valid_and_not_has_been_sent & mm__done_load_en;
  assign tmp4 = {tmp4__2, ____state_3};
  assign tmp8 = {add_667, ____state_2[1:0]};
  assign tmp18 = p3_slt_687 ? tmp17 : tmp3;
  assign mm__go_load_en = mm__go_vld & mm__go_valid_load_en;
  assign mm__mem0__read_resp_load_en = mm__mem0__read_resp_vld & mm__mem0__read_resp_valid_load_en;
  assign mm__mem1__read_resp_load_en = mm__mem1__read_resp_vld & mm__mem1__read_resp_valid_load_en;
  assign mm__mem2__write_resp_load_en = mm__mem2__write_resp_vld & mm__mem2__write_resp_valid_load_en;
  assign or_1221 = ~p0_stage_done | ____state_0__at_most_one_next_value | rst;
  assign or_1223 = ~p0_stage_done | ____state_1__at_most_one_next_value | rst;
  assign or_1225 = ~p0_stage_done | ____state_2__at_most_one_next_value | rst;
  assign or_1227 = ~p0_stage_done | ____state_3__at_most_one_next_value | rst;
  assign or_679 = ____state_3[0] | ____state_3[1];
  assign tmp21 = {add_699, ____state_2[1:0]};
  assign and_712 = tmp20 & slt_688;
  assign one_hot_sel_1040 = tmp2 & {32{concat_1039[0]}} | tmp17 & {32{concat_1039[1]}} | tmp2 & {32{concat_1039[2]}};
  assign or_1041 = and_1035 | and_1036 | and_1037;
  assign one_hot_sel_1047 = add_682 & {32{concat_1046[0]}} | tmp2 & {32{concat_1046[1]}};
  assign or_1048 = and_1043 | and_1044;
  assign one_hot_sel_1054 = add_681 & {32{concat_1053[0]}} | tmp2 & {32{concat_1053[1]}};
  assign or_1055 = and_1050 | and_1051;
  assign tmp32 = tmp1 | ____state_4 & nand_690;
  assign one_hot_sel_1061 = unexpand_for_next_value_158_3_case_1 & {2{concat_1060[0]}} | unexpand_for_next_value_158_3_case_0 & {2{concat_1060[1]}};
  assign or_1062 = and_1058 | and_1059;
  assign __mm__mem0__read_req_not_stage_load = ~__mm__mem0__read_req_valid_and_all_active_outputs_ready;
  assign __mm__mem0__read_req_has_been_sent_reg_load_en = __mm__mem0__read_req_valid_and_ready_txfr | __mm__mem0__read_req_valid_and_all_active_outputs_ready;
  assign __mm__mem1__read_req_has_been_sent_reg_load_en = __mm__mem1__read_req_valid_and_ready_txfr | __mm__mem0__read_req_valid_and_all_active_outputs_ready;
  assign __mm__mem2__write_req_not_stage_load = ~__mm__mem2__write_req_valid_and_all_active_outputs_ready;
  assign __mm__mem2__write_req_has_been_sent_reg_load_en = __mm__mem2__write_req_valid_and_ready_txfr | __mm__mem2__write_req_valid_and_all_active_outputs_ready;
  assign __mm__done_not_stage_load = ~__mm__done_valid_and_all_active_outputs_ready;
  assign __mm__done_has_been_sent_reg_load_en = __mm__done_valid_and_ready_txfr | __mm__done_valid_and_all_active_outputs_ready;
  assign tmp5 = {tmp4};
  assign tmp9 = {tmp8};
  assign tmp23 = {p3_tmp21, tmp18};
  assign __mm__done_buf = 1'h1;
  always_ff @ (posedge clk) begin
    if (rst) begin
      ____state_2 <= 32'h0000_0000;
      ____state_1 <= 32'h0000_0000;
      ____state_3 <= 2'h0;
      ____state_4 <= 1'h0;
      p0_or_679 <= 1'h0;
      p0_slt_687 <= 1'h0;
      p0_tmp21 <= 4'h0;
      p0_and_712 <= 1'h0;
      p0_tmp27 <= 1'h0;
      p0_and_701 <= 1'h0;
      p0_and_702 <= 1'h0;
      p1_or_679 <= 1'h0;
      p1_slt_687 <= 1'h0;
      p1_tmp21 <= 4'h0;
      p1_and_712 <= 1'h0;
      p1_tmp27 <= 1'h0;
      p1_and_701 <= 1'h0;
      p1_and_702 <= 1'h0;
      p2_or_679 <= 1'h0;
      p2_slt_687 <= 1'h0;
      p2_tmp21 <= 4'h0;
      p2_and_712 <= 1'h0;
      p2_tmp27 <= 1'h0;
      p2_and_701 <= 1'h0;
      p2_and_702 <= 1'h0;
      p3_or_679 <= 1'h0;
      p3_slt_687 <= 1'h0;
      p3_tmp21 <= 4'h0;
      p3_and_712 <= 1'h0;
      p3_tmp27 <= 1'h0;
      p3_and_701 <= 1'h0;
      p3_and_702 <= 1'h0;
      ____state_0 <= 32'h0000_0000;
      p4_and_712 <= 1'h0;
      p4_tmp27 <= 1'h0;
      p5_and_712 <= 1'h0;
      p5_tmp27 <= 1'h0;
      p6_and_712 <= 1'h0;
      p6_tmp27 <= 1'h0;
      p7_and_712 <= 1'h0;
      p7_tmp27 <= 1'h0;
      p0_valid <= 1'h0;
      p1_valid <= 1'h0;
      p2_valid <= 1'h0;
      p3_valid <= 1'h0;
      p4_valid <= 1'h0;
      p5_valid <= 1'h0;
      p6_valid <= 1'h0;
      p7_valid <= 1'h0;
      __mm__mem0__read_req_has_been_sent_reg <= 1'h0;
      __mm__mem1__read_req_has_been_sent_reg <= 1'h0;
      __mm__mem2__write_req_has_been_sent_reg <= 1'h0;
      __mm__done_has_been_sent_reg <= 1'h0;
      __mm__go_reg <= 1'h0;
      __mm__go_valid_reg <= 1'h0;
      __mm__mem0__read_resp_reg <= __mm__mem0__read_resp_reg_init;
      __mm__mem0__read_resp_valid_reg <= 1'h0;
      __mm__mem1__read_resp_reg <= __mm__mem1__read_resp_reg_init;
      __mm__mem1__read_resp_valid_reg <= 1'h0;
      __mm__mem2__write_resp_valid_reg <= 1'h0;
      __mm__mem0__read_req_reg <= __mm__mem0__read_req_reg_init;
      __mm__mem0__read_req_valid_reg <= 1'h0;
      __mm__mem1__read_req_reg <= __mm__mem1__read_req_reg_init;
      __mm__mem1__read_req_valid_reg <= 1'h0;
      __mm__mem2__write_req_reg <= __mm__mem2__write_req_reg_init;
      __mm__mem2__write_req_valid_reg <= 1'h0;
      __mm__done_reg <= 1'h0;
      __mm__done_valid_reg <= 1'h0;
    end else begin
      ____state_2 <= or_1055 ? one_hot_sel_1054 : ____state_2;
      ____state_1 <= or_1048 ? one_hot_sel_1047 : ____state_1;
      ____state_3 <= or_1062 ? one_hot_sel_1061 : ____state_3;
      ____state_4 <= p0_data_enable ? tmp32 : ____state_4;
      p0_or_679 <= p0_data_enable ? or_679 : p0_or_679;
      p0_slt_687 <= p0_data_enable ? slt_687 : p0_slt_687;
      p0_tmp21 <= p0_data_enable ? tmp21 : p0_tmp21;
      p0_and_712 <= p0_data_enable ? and_712 : p0_and_712;
      p0_tmp27 <= p0_data_enable ? tmp27 : p0_tmp27;
      p0_and_701 <= p0_data_enable ? and_701 : p0_and_701;
      p0_and_702 <= p0_data_enable ? and_702 : p0_and_702;
      p1_or_679 <= p1_data_enable ? p0_or_679 : p1_or_679;
      p1_slt_687 <= p1_data_enable ? p0_slt_687 : p1_slt_687;
      p1_tmp21 <= p1_data_enable ? p0_tmp21 : p1_tmp21;
      p1_and_712 <= p1_data_enable ? p0_and_712 : p1_and_712;
      p1_tmp27 <= p1_data_enable ? p0_tmp27 : p1_tmp27;
      p1_and_701 <= p1_data_enable ? p0_and_701 : p1_and_701;
      p1_and_702 <= p1_data_enable ? p0_and_702 : p1_and_702;
      p2_or_679 <= p2_data_enable ? p1_or_679 : p2_or_679;
      p2_slt_687 <= p2_data_enable ? p1_slt_687 : p2_slt_687;
      p2_tmp21 <= p2_data_enable ? p1_tmp21 : p2_tmp21;
      p2_and_712 <= p2_data_enable ? p1_and_712 : p2_and_712;
      p2_tmp27 <= p2_data_enable ? p1_tmp27 : p2_tmp27;
      p2_and_701 <= p2_data_enable ? p1_and_701 : p2_and_701;
      p2_and_702 <= p2_data_enable ? p1_and_702 : p2_and_702;
      p3_or_679 <= p3_data_enable ? p2_or_679 : p3_or_679;
      p3_slt_687 <= p3_data_enable ? p2_slt_687 : p3_slt_687;
      p3_tmp21 <= p3_data_enable ? p2_tmp21 : p3_tmp21;
      p3_and_712 <= p3_data_enable ? p2_and_712 : p3_and_712;
      p3_tmp27 <= p3_data_enable ? p2_tmp27 : p3_tmp27;
      p3_and_701 <= p3_data_enable ? p2_and_701 : p3_and_701;
      p3_and_702 <= p3_data_enable ? p2_and_702 : p3_and_702;
      ____state_0 <= or_1041 ? one_hot_sel_1040 : ____state_0;
      p4_and_712 <= p4_data_enable ? p3_and_712 : p4_and_712;
      p4_tmp27 <= p4_data_enable ? p3_tmp27 : p4_tmp27;
      p5_and_712 <= p5_data_enable ? p4_and_712 : p5_and_712;
      p5_tmp27 <= p5_data_enable ? p4_tmp27 : p5_tmp27;
      p6_and_712 <= p6_data_enable ? p5_and_712 : p6_and_712;
      p6_tmp27 <= p6_data_enable ? p5_tmp27 : p6_tmp27;
      p7_and_712 <= p7_data_enable ? p6_and_712 : p7_and_712;
      p7_tmp27 <= p7_data_enable ? p6_tmp27 : p7_tmp27;
      p0_valid <= p0_enable ? p0_stage_done : p0_valid;
      p1_valid <= p1_enable ? p0_valid : p1_valid;
      p2_valid <= p2_enable ? p1_valid : p2_valid;
      p3_valid <= p3_enable ? p2_valid : p3_valid;
      p4_valid <= p4_enable ? p4_stage_done : p4_valid;
      p5_valid <= p5_enable ? p4_valid : p5_valid;
      p6_valid <= p6_enable ? p5_valid : p6_valid;
      p7_valid <= p7_enable ? p6_valid : p7_valid;
      __mm__mem0__read_req_has_been_sent_reg <= __mm__mem0__read_req_has_been_sent_reg_load_en ? __mm__mem0__read_req_not_stage_load : __mm__mem0__read_req_has_been_sent_reg;
      __mm__mem1__read_req_has_been_sent_reg <= __mm__mem1__read_req_has_been_sent_reg_load_en ? __mm__mem0__read_req_not_stage_load : __mm__mem1__read_req_has_been_sent_reg;
      __mm__mem2__write_req_has_been_sent_reg <= __mm__mem2__write_req_has_been_sent_reg_load_en ? __mm__mem2__write_req_not_stage_load : __mm__mem2__write_req_has_been_sent_reg;
      __mm__done_has_been_sent_reg <= __mm__done_has_been_sent_reg_load_en ? __mm__done_not_stage_load : __mm__done_has_been_sent_reg;
      __mm__go_reg <= mm__go_load_en ? mm__go : __mm__go_reg;
      __mm__go_valid_reg <= mm__go_valid_load_en ? mm__go_vld : __mm__go_valid_reg;
      __mm__mem0__read_resp_reg <= mm__mem0__read_resp_load_en ? mm__mem0__read_resp : __mm__mem0__read_resp_reg;
      __mm__mem0__read_resp_valid_reg <= mm__mem0__read_resp_valid_load_en ? mm__mem0__read_resp_vld : __mm__mem0__read_resp_valid_reg;
      __mm__mem1__read_resp_reg <= mm__mem1__read_resp_load_en ? mm__mem1__read_resp : __mm__mem1__read_resp_reg;
      __mm__mem1__read_resp_valid_reg <= mm__mem1__read_resp_valid_load_en ? mm__mem1__read_resp_vld : __mm__mem1__read_resp_valid_reg;
      __mm__mem2__write_resp_valid_reg <= mm__mem2__write_resp_valid_load_en ? mm__mem2__write_resp_vld : __mm__mem2__write_resp_valid_reg;
      __mm__mem0__read_req_reg <= mm__mem0__read_req_load_en ? tmp5 : __mm__mem0__read_req_reg;
      __mm__mem0__read_req_valid_reg <= mm__mem0__read_req_valid_load_en ? __mm__mem0__read_req_valid_and_not_has_been_sent : __mm__mem0__read_req_valid_reg;
      __mm__mem1__read_req_reg <= mm__mem1__read_req_load_en ? tmp9 : __mm__mem1__read_req_reg;
      __mm__mem1__read_req_valid_reg <= mm__mem1__read_req_valid_load_en ? __mm__mem1__read_req_valid_and_not_has_been_sent : __mm__mem1__read_req_valid_reg;
      __mm__mem2__write_req_reg <= mm__mem2__write_req_load_en ? tmp23 : __mm__mem2__write_req_reg;
      __mm__mem2__write_req_valid_reg <= mm__mem2__write_req_valid_load_en ? __mm__mem2__write_req_valid_and_not_has_been_sent : __mm__mem2__write_req_valid_reg;
      __mm__done_reg <= mm__done_load_en ? __mm__done_buf : __mm__done_reg;
      __mm__done_valid_reg <= mm__done_valid_load_en ? __mm__done_valid_and_not_has_been_sent : __mm__done_valid_reg;
    end
  end
  assign mm__done = __mm__done_reg;
  assign mm__done_vld = __mm__done_valid_reg;
  assign mm__go_rdy = mm__go_load_en;
  assign mm__mem0__read_req = __mm__mem0__read_req_reg;
  assign mm__mem0__read_req_vld = __mm__mem0__read_req_valid_reg;
  assign mm__mem0__read_resp_rdy = mm__mem0__read_resp_load_en;
  assign mm__mem1__read_req = __mm__mem1__read_req_reg;
  assign mm__mem1__read_req_vld = __mm__mem1__read_req_valid_reg;
  assign mm__mem1__read_resp_rdy = mm__mem1__read_resp_load_en;
  assign mm__mem2__write_req = __mm__mem2__write_req_reg;
  assign mm__mem2__write_req_vld = __mm__mem2__write_req_valid_reg;
  assign mm__mem2__write_resp_rdy = mm__mem2__write_resp_load_en;
  `ifdef ASSERT_ON
  ____state_0__at_most_one_next_value_assert: assert property (@(posedge clk) disable iff ($sampled(rst !== 1'h0 || $isunknown(or_1221))) or_1221) else $fatal(0, "More than one next_value fired for state element: __state_0");
  ____state_1__at_most_one_next_value_assert: assert property (@(posedge clk) disable iff ($sampled(rst !== 1'h0 || $isunknown(or_1223))) or_1223) else $fatal(0, "More than one next_value fired for state element: __state_1");
  ____state_2__at_most_one_next_value_assert: assert property (@(posedge clk) disable iff ($sampled(rst !== 1'h0 || $isunknown(or_1225))) or_1225) else $fatal(0, "More than one next_value fired for state element: __state_2");
  ____state_3__at_most_one_next_value_assert: assert property (@(posedge clk) disable iff ($sampled(rst !== 1'h0 || $isunknown(or_1227))) or_1227) else $fatal(0, "More than one next_value fired for state element: __state_3");
  `endif  // ASSERT_ON
endmodule
